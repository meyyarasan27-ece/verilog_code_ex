`timescale 1ns / 1ps
module mux16_1_tb();
reg i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15 ;
reg s0,s1,s2,s3 ;
wire y ;

mux16_1 dut (
  .i0(i0), .i1(i1), .i2(i2), .i3(i3),
  .i4(i4), .i5(i5), .i6(i6), .i7(i7),
  .i8(i8), .i9(i9), .i10(i10), .i11(i11),
  .i12(i12), .i13(i13), .i14(i14), .i15(i15),
  .s0(s0), .s1(s1), .s2(s2), .s3(s3),
  .y(y)
);

initial begin
$monitor(" time = %t || i0 = %b || i1  = %b|| i2 = %b || i3 = %b || i4 = %b || i5 = %b || i6 = %b || i7 = %b || i8 = %b || i9 = %b || i10 = %b || i11 = %b || i12 = %b || i13 = %b || i14  = %b || i15 = %b || s3 = %b || s2 = %b || s1 = %b || s0 = %b || y = %b ",$time ,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15 ,s3,s2,s1,s0,y);

i0 = 1'b0 ;i1 = 1'b1 ;i2 = 1'b0 ;i3 = 1'b1 ;
i4 = 1'b0; i5 = 1'b1 ;i6 = 1'b1 ;i7 = 1'b0 ;
i8 = 1'b1 ;i9 = 1'b0 ;i10 = 1'b1 ;i11 = 1'b1 ;
i12 = 1'b1 ;i13 = 1'b0 ;i14 = 1'b1 ;i15  = 1'b0 ;


 s0 = 1'b0 ;s1 = 1'b0 ; s2 =1'b0 ; s3 = 1'b0 ; #10 ;
s0 = 1'b0 ;s1 = 1'b0 ; s2 = 1'b0 ; s3 = 1'b1 ; #10;
s0 = 1'b0 ;s1 = 1'b0 ; s2 = 1'b1 ; s3 = 1'b0 ; #10;
s0 = 1'b0 ;s1 = 1'b0 ; s2 = 1'b1 ; s3 = 1'b1 ; #10;
s0 = 1'b0 ;s1 = 1'b1 ; s2 = 1'b0 ; s3 = 1'b0 ; #10;
s0 = 1'b0 ;s1 = 1'b1 ; s2 = 1'b0 ; s3 = 1'b1 ; #10;
s0 = 1'b0 ;s1 = 1'b1 ; s2 = 1'b1 ; s3 = 1'b0 ; #10;
s0 = 1'b0 ;s1 = 1'b1 ; s2 = 1'b1 ; s3 = 1'b1 ; #10;
s0 = 1'b1 ;s1 = 1'b0 ; s2 = 1'b0 ; s3 = 1'b0 ; #10;
s0 = 1'b1 ;s1 = 1'b0 ; s2 = 1'b0 ; s3 = 1'b1 ; #10;
s0 = 1'b1 ;s1 = 1'b0 ; s2 = 1'b1 ; s3 = 1'b0 ; #10;
s0 = 1'b1 ;s1 = 1'b0 ; s2 = 1'b1 ; s3 = 1'b1 ; #10;
s0 = 1'b1 ;s1 = 1'b1 ; s2 = 1'b0 ; s3 = 1'b0 ; #10;
s0 = 1'b1 ;s1 = 1'b1 ; s2 = 1'b0 ; s3 = 1'b1 ; #10;
s0 = 1'b1 ;s1 = 1'b1 ; s2 = 1'b1 ; s3 = 1'b0 ; #10;
s0 = 1'b1 ;s1 = 1'b1 ; s2 = 1'b1 ; s3 = 1'b1 ; #10;

$finish;
end
endmodule
